// Top module of USI

//test branch