// Top level testbench for USI
module top_tb();

endmodule