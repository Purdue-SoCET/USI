// Top module of USI