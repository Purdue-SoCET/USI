module reg_map(
    input logic CLK,
    input logic nRST
)

endmodule