// Top level testbench for USI