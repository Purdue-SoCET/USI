module reg_map_tb();

endmodule